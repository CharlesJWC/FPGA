//`include "Memory.v"

module tb_MIPS;

reg CLK;
wire CS, WE;

parameter N = 10;
reg [31:0] expected[N:1];

wire[31:0] Address, Address_MUX, Mem_Bus_Wire;
reg[31:0] AddressTB;
wire WE_MUX, CS_MUX;
reg init, rst, WE_TB, CS_TB;

integer i;

MIPS CPU(CLK,rst, CS, WE, Address, Mem_Bus_Wire);
Memory MEM(CS_MUX, WE_MUX, CLK, Address_MUX, Mem_Bus_Wire);

assign Address_MUX = (init)? AddressTB: Address;
assign WE_MUX = (init)? WE_TB : WE;
assign CS_MUX = (init)? CS_TB : CS;

always #10 CLK = ~CLK;

initial 
begin
	expected[1] = 32'h00000006;	// 6
	expected[2] = 32'h00000012;	// 18
	expected[3] = 32'h00000018;	// 24
	expected[4] = 32'h0000000C;	// 12
	expected[5] = 32'h00000002;	// 2
	expected[6] = 32'h00000016;	// 22
	expected[7] = 32'h00000001;	// 1
	expected[8] = 32'h00000120;	// 288
	expected[9] = 32'h00000003;	// 3
	expected[10] = 32'h00412022;// 5th Instruction
	CLK = 0;
end

always 
begin

	rst = 1;
	@(posedge CLK);
	init <=1; CS_TB<=1; WE_TB<=1;
	@(posedge CLK);
	CS_TB<=0; WE_TB<=0; init <=0;
	@(posedge CLK);
	rst <= 0;
	for(i = 1; i <= N; i = i+1)
	begin
		@(posedge WE);
		@(negedge CLK);
		if(Mem_Bus_Wire != expected[i])
			$display("result Mismatch!\n got : %d\t expect : %d",Mem_Bus_Wire,expected[i]);
	end
	$display("Testing Finished!");
	$stop;
end
endmodule 