module tb_upcounter_4bits;

reg t_clk;
reg t_rst;
reg t_up;
wire [3:0] t_q;


upcounter_4bits t_upcounter_4bits
(
	.clk(t_clk),
	.rst(t_rst),
	.up(t_up),
	.q(t_q)
);


initial
begin
	t_clk = 1'b1;
	t_rst = 1'b1;
	t_up = 1'b0;
end

always
begin
	#3 t_clk = ~t_clk;
end

initial
begin
	#3  t_rst = 1'b0; t_up = 1'b1;
	#30 t_up = 1'b0;
	#9  t_up = 1'b1;
	#15 t_rst = 1'b1;
	#18 t_rst = 1'b0;
	#24 t_rst = 1'b1;
	#3  t_rst = 1'b0;
end

endmodule
	
	
	

	