module MIPS
(
	input clk,
	input [15:0] Instr,
	output current_state
);





