module mux_4x1 (in0, in1, in2, in3, select, out);

input in0, in1, in2, in3;
input [1:0] select;
output out;

assign out = select[1] ? (select[0] ? in3 : in2) : (select[0] ? in1 : in0);


endmodule
