module tb_deconder_2x4;
// 2x4 ���ڴ� ��� �ùķ��̼��� ���� �׽�Ʈ��ġ ��� ����

reg [1:0] t_in; // 2bits �Է� ��ȣ ��Ʈ ����
reg t_enable; // EN ��ȣ �Է� ��Ʈ ����
// �� �Է� ��ȣ�� ��ȭ��ų �� �ֵ��� reg������ ���� 
wire [3:0] t_out; // 4bits ��� ��Ʈ ����
// ���ڴ� ����� ��� ���� �޾� ��¸� �ϸ� �ǹǷ� wire������ ����

decoder_2x4 t_decoder_2x4 // 2x4 ���ڴ� ��� ��ü ����
(
	// ����� �� ����� ��Ʈ�� �ù����̼� ��Ʈ�� �̸��� ���� ����
	.in(t_in),
	.enable(t_enable),
	.out(t_out)
);

initial // t = 0�� �� ��� �Է°� �ʱ�ȭ
begin
	t_in = 2'd0;		//00
	t_enable = 1'b0;	//1(high)
end

always	// t = 0 �� ������ 40ns���� EN��ȣ ��ȭ(Toggle)
begin
	#40 t_enable = ~t_enable;
end

always // t = 0 �� ������ 10ns���� �Է� ��ȣ ��ȭ
begin 
#0	t_in = 2'd0; #10;	//00 -- EN��ȣ High�� ��
// �Է� ��ȣ �ʱ�ȭ�� Ȯ���ϰ� �Ϸ�� ���� �Է� ��ȣ�� �ֱ� ���Ͽ� #0 �߰�
	t_in = 2'd1; #10;	//01
	t_in = 2'd2; #10;	//10
	t_in = 2'd3; #10;	//11
	t_in = 2'd0; #10;	//00 -- EN��ȣ Low�� ��
	t_in = 2'd1; #10;	//01
	t_in = 2'd2; #10;	//10
	t_in = 2'd3; #10;	//11
end

endmodule // 2x4 ���ڴ� �׽�Ʈ��ġ ��� ��� �Ϸ�