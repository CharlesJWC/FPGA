module fullAdder
(
	sum,
	c_out,
	a,
	b,
	c_in
);

input a;
input b;
input c_in;
output sum;
output c_out;

wire s1, s2, c1;

xor(s1, a, b);
and(c1, a, b);
xor(sum, s1, c_in);
and(s2, s1, c_in);
or(c_out, s2, c1);

endmodule


